module sd_read(
    output reg sd_clk,
    inout sd_dat0,
    inout sd_cmd
);

// TODO
// https://web.archive.org/web/20200725013613/http://wiki.seabright.co.nz/wiki/SdCardProtocol.html

endmodule
